uvm _reg  TOTAL_CREDIT  // Total power credit for flash active control (BLG_Rbase + 0x00), offset = (BLG_Rbase + 0x00)
uvm _reg  CW_SIZE  // Code Word Size (BLG_Rbase + 0x04), offset = (BLG_Rbase + 0x04)
uvm _reg  CW_ZERO  // Code Word zero bit limit (BLG_Rbase + 0x08), offset = (BLG_Rbase + 0x08)
uvm _reg  C0_REMAP  // Remap Channel 0 Address to other channel (BLG_Rbase + 0x0C), offset = (BLG_Rbase + 0x0C)
uvm _reg  Spare_Reg  // Spare register (BLG_Rbase + 0x10), offset = (BLG_Rbase + 0x10)
uvm _reg  Sys_freq  // System Frequency (BLG_Rbase + 0x14), offset = (BLG_Rbase + 0x14)
uvm _reg  FPH_Pow_itv  // Re-request Power Interval (BLG_Rbase + 0x18), offset = (BLG_Rbase + 0x18)
uvm _reg  FPH_CE_IDLE  // FPH CE Idle value (BLG_Rbase + 0x1C), offset = (BLG_Rbase + 0x1C)
uvm _reg  FPH_INT_SRC  // FPH Interrupt source (BLG_Rbase + 0x20), offset = (BLG_Rbase + 0x20)
uvm _reg  FPH_INT_RAW  // FPH Interrupt Raw Data (BLG_Rbase + 0x24), offset = (BLG_Rbase + 0x24)
uvm _reg  FPH_INT_EN  // FPH Interrupt Raw Data (GLB_Rbase + 0x28), offset = (GLB_Rbase + 0x28)
uvm _reg  FPH_INT_DBG  // FPH Interrupt Debug (GLB_Rbase + 0x2C), offset = (GLB_Rbase + 0x2C)
uvm _reg  MTC_DBG_CFG  // MTC Debug Config (GLB_Rbase + 0x30), offset = (GLB_Rbase + 0x30)
uvm _reg  MTC_DBG_BADDR  // MTC Debug  Base Addr (GLB_Rbase + 0x34), offset = (GLB_Rbase + 0x34)
uvm _reg  MTC_DBG_WPTR  // MTC Debug  Write Point (GLB_Rbase + 0x38), offset = (GLB_Rbase + 0x38)
uvm _reg  MTC_DBG_WPTR  // FPH Debug Fake ADT (GLB_Rbase + 0x3C), offset = (GLB_Rbase + 0x3C)
uvm _reg  MTC_DBG_SQ  // MTC Debug SQ_0~7  (GLB_Rbase + 0x40 ~ 0x5C), offset = (GLB_Rbase + 0x40)
uvm _reg  MTC_DBG_SQ_Trig  // MTC Debug SQ_Trigger + 0x60, offset = (none + none)
uvm _reg  FPH_DBG_Fake_ADM_CWL  // FPH Debug Fake ADM CW Value L (GLB_Rbase + 0x70), offset = (GLB_Rbase + 0x70)
uvm _reg  FPH_DBG_Fake_ADM_CWH  // FPH Debug Fake ADM CW Value H (GLB_Rbase + 0x74), offset = (GLB_Rbase + 0x74)
uvm _reg  FPH_IO_RBN  // FPH IP Rdy Busy  (GLB_Rbase + 0x78), offset = (GLB_Rbase + 0x78)
uvm _reg  FPH_PWR_LOSS  // FPH Power Loss Flag  (GLB_Rbase + 0x7C), offset = (GLB_Rbase + 0x7C)
uvm _reg  FPH_CH_LRdata  // FPH Channel Last Read data   (GLB_Rbase + 0x80~0x9C), offset = (GLB_Rbase + 0x80~0x9C)
uvm _reg  FPH_ADM_IF_Watch  // FPH ADM IF Watch Signal   (GLB_Rbase + 0xA0~0xBC), offset = (GLB_Rbase + 0xA0~0xBC)
uvm _reg  FPH_CH_STOP  // FPH Channel Stop   (GLB_Rbase + 0xD0), offset = (GLB_Rbase + 0xD0)
uvm _reg  FPH_CH_MTC_Exec  // FPH Channel MTC Exec   (GLB_Rbase + 0xD4), offset = (GLB_Rbase + 0xD4)
uvm _reg  FPH_CH_MTC_Exec  // FPH Select Debug MTC Channel   (GLB_Rbase + 0xD8), offset = (GLB_Rbase + 0xD8)
uvm _reg  FPH_Dbg_Curr_MTC  // FPH Debug Current Exec MTC   (GLB_Rbase + 0xE0~0xFC), offset = (GLB_Rbase + 0xE0~0xFC)
uvm _reg  FPH_Time_First_Pol  //  FPH Timer First Polling   (GLB_Rbase + 0x100 ~0x10C), offset = (GLB_Rbase + 0x100)
uvm _reg  FPH_Timeout_CFG  // FPH Timeout Config   (GLB_Rbase + 0x110 ~0x11C), offset = (GLB_Rbase + 0x110)
uvm _reg  FPH_Time_Pol_Interval  // FPH Timer Polling Interval   (GLB_Rbase + 0x120), offset = (GLB_Rbase + 0x120)
uvm _reg  FPH_Time_Pol_Interval  // FPH Write Page Dummy Enable  (GLB_Rbase + 0x130), offset = (GLB_Rbase + 0x130)
uvm _reg  FPH_Wpage_Dummy_Length  // FPH Write Page Dummy Lenght  (GLB_Rbase + 0x134), offset = (GLB_Rbase + 0x134)
uvm _reg  FPH_High_QNUM  // FPH High Priority Queue Number  (GLB_Rbase + 0x500~0x51C), offset = (GLB_Rbase + 0x500~0x51C)

uvm _reg  PIO_ENABLE  // Set up the FPH PIO mode, offset = (none + none)
uvm _reg  PIO_TAG  // Trigger the FPH send the TAG to ADM, offset = (Chx_Rbase + 0x04)
uvm _reg  PIO_BUF_ST  // PIO buffer status, offset = (Chx_Rbase + 0x08)
uvm _reg  MTC_CE_MAP_CE_0  // MTC Queue Mapping CE 0, offset = (Chx_Rbase + 0x10)
uvm _reg  MTC_CE_MAP_CE_1  // MTC Queue Mapping CE_1, offset = (Chx_Rbase + 0x14)
uvm _reg  MTC_CE_MAP_CE_2  // MTC Queue Mapping CE_2, offset = (Chx_Rbase + 0x18)
uvm _reg  MTC_CE_MAP_CE_3  // MTC Queue Mapping CE_3, offset = (Chx_Rbase + 0x1C)
uvm _reg  MTC_CE_MAP_CE_4  // MTC Queue Mapping CE_4, offset = (Chx_Rbase + 0x20)
uvm _reg  MTC_CE_MAP_CE_5  // MTC Queue Mapping CE_5, offset = (Chx_Rbase + 0x24)
uvm _reg  MTC_CE_MAP_CE_6  // MTC Queue Mapping CE_6, offset = (Chx_Rbase + 0x28)
uvm _reg  MTC_CE_MAP_CE_7  // MTC Queue Mapping CE_7, offset = (Chx_Rbase + 0x2C)
uvm _reg  MTC_CE_MAP_CE_8  // MTC Queue Mapping CE_8, offset = (Chx_Rbase + 0x30)
uvm _reg  MTC_CE_MAP_CE_9  // MTC Queue Mapping CE_9, offset = (Chx_Rbase + 0x34)
uvm _reg  MTC_CE_MAP_CE_10  // MTC Queue Mapping CE_10, offset = (Chx_Rbase + 0x38)
uvm _reg  MTC_CE_MAP_CE_11  // MTC Queue Mapping CE_11, offset = (Chx_Rbase + 0x3C)
uvm _reg  MTC_CE_MAP_CE_10  // MTC Queue Mapping CE_10, offset = (Chx_Rbase + 0x38)
uvm _reg  MTC_CE_MAP_CE_31  // MTC Queue Mapping CE_31, offset = (Chx_Rbase + 0x8C)
uvm _reg  MTC_FPHY_TIME  // MTC FPHY TIME Setting, offset = (Chx_Rbase + 0x90)
uvm _reg  MTC_FPHY_MODE  // MTC FPHY mode Setting, offset = (Chx_Rbase + 0x94)
uvm _reg  NO_MTC_HOLD  // Normal queue MTC Hold, offset = (Chx_Rbase + 0x98)
uvm _reg  HQ_MTC_HOLD  // High priority Queue MTC Hold, offset = (Chx_Rbase + 0x9C)
uvm _reg  NO_MTC_STEP  // Normal queue MTC step, offset = (Chx_Rbase + 0xA4)
uvm _reg  HQ_MTC_STEP  // High priority Queue MTC Step, offset = (Chx_Rbase + 0xA8)
uvm _reg  FCU_Rdata  // FCU Rdata Register, offset = (none + none)
uvm _reg  FCU_CState  // FCU Current State, offset = (none + none)
uvm _reg  FCU_CFCUAddr  // FCU Current FCU Addr, offset = (none + none)
uvm _reg  FCU_Mode_EN  // FCU Mode Enable, offset = (none + none)
uvm _reg  FCU_Cmd  // FCU Command, offset = (none + none)
uvm _reg  FCU_CK_Switch  // FCU Clock Switch, offset = (Chx_Rbase + 0xC4)

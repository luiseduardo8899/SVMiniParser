

typedef struct packed {	 

    bit [95:32] PPA;
    bit [31:24] IDX;
    bit [23:20] SPLIT_ID;
    bit [15:0] CTAG;
    
} to_MEC_PPA_s;

